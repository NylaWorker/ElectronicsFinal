`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:54:48 11/08/2017 
// Design Name: 
// Module Name:    pmodExploration 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pmodExploration(a,b);
	(*LOC = "A8" *) input  a;
	(*LOC = "N10" *) output b;
	assign b = a; 


endmodule
